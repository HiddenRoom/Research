include "../instructionDecode.v"

module test_instructionDecode.v;


endmodule