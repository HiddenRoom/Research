`ifndef __REGFILE__
`define __REGFILE__

module regFile
(
  input [4:0]     read0,
  input [4:0]     read1,
  input [4:0]     read2,
  input [4:0]     read3,
);


module

`endif
