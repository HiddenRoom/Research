include "../alu.v"

module test_alu.v;


endmodule