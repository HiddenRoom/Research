`ifndef __PRIORITYROUTER__
`define __PRIORITYROUTER__

module
(
  // take in input val and version num and read input with version num and
  // output the nearest version inside with a version num less than input
  // version num 
);

endmodule

`endif
