include "../priorityRouter.v"

module test_priorityRouter.v;


endmodule